/* verilator lint_off UNUSEDPARAM */
localparam MEMW_BYTE = 2'b00;
localparam MEMW_HALF = 2'b01;
localparam MEMW_WORD = 2'b10;
/* verilator lint_on UNUSEDPARAM */
